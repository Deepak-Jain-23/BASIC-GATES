// Code your design here
module basicgates(a,b,y1,y2,y3,y4,y5,y6,y7);
  input  a;
  input  b;
  output  y1,y2,y3,y4,y5,y6,y7;
  and(y1,a,b);
or(y2,a,b);
not(y3,a);
nand(y4,a,b);
nor(y5,a,b);
xor(y6,a,b);
xnor(y7,a,b);
endmodule